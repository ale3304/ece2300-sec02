//========================================================================
// PairTripleDetector
//========================================================================

//test comment 

module PairTripleDetector
(
  input  wire in0,
  input  wire in1,
  input  wire in2,
  output wire out
);
  // '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''
  // Discussion Section Task
  // '''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''''
  // Implement a pair/triple detector using explicit gate-level modeling.
assign out = (~in0 && in1 && in2) || (in0 && ~in1 && in2) || (in0 && in1 && ~in2) || (in0 && in1 && in2);

endmodule

